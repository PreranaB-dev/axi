//================================================================
//---------AXI_DEFINES-------------
// Description : This file has all the defines used inside the
//               rtl main code. Define all parameters here.
// Warning     : No gurantee. Use at your own risk.
//================================================================

//
`define DATA_BITS  32
`define ADDR_BITS  32
`define LEN_BITS   1
`define SIZE_BITS  1

