//---------------------------------
//---------AXI_DEFINES-------------
//---------------------------------
//---12july2020-------------

`define DATA_BITS 
`define ADDR_BITS
`define LEN_BITS
`define SIZE_BITS

